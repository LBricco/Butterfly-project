--**********************************************************************************
--* Micro ROM per la microprogrammazione della control unit
--* Ogni riga è costituita da 36 bit
--* Bit 35-7: segnali di controllo che governano il funzioanmento del circuito
--* Bit 6-2: jump address
--* Bit 1-0: condition code
--**********************************************************************************

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity uROM_butterfly is
    port (
        ADDR : in integer range 0 to 19;
        CELL : out std_logic_vector(42 downto 0)
    );
end entity uROM_butterfly;

architecture structure of uROM_butterfly is

    type rom is array (0 to 19) of std_logic_vector(42 downto 0);
    constant micro_rom : rom := (
        "1111110000100000000000000000000000100000000",
        "0000000000100000000000100000000000000000000",
        "0000000000101000000000100000000000000000000",
        "0000000000111000100000100000000000000000000",
        "0000000000110000100000110000000000000000000",
        "0010001000000100100000010000001101100000000",
        "1111110000010011100100001000000000000000000",
        "0000000000100001100010100000000000000000000",
        "0000000000101010110001100110000000000000000",
        "0000100010111001101000100011000000000000000",
        "0000110011110000100000110001000000000000000",
        "0010101100000100100000010000000000000000000",
        "0000000000010011100100001000100110110111010",
        "0000000000010011100100001000000000000000000",
        "0000000000000001100010000000000000000000000",
        "0000000000000010110001000110000000000000000",
        "0000100010000001001000000011000000000000000",
        "0000110011000000000000000001000000000000000",
        "0000100100000000000000000000000000000000000",
        "0000000000000000000000000000100000010000000"

    );

begin

    CELL <= micro_rom(ADDR);

end architecture structure;